/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   framebuffer.cdl
 * @brief  Framebuffer module with separate display and video sides
 *
 * CDL implementation of a module that takes SRAM writes into a
 * framebuffer, and includes a mapping to a dual-port SRAM (write on
 * one side, read on the other), where the video side drives out
 * vsync, hsync, data enable and pixel data.
 *
 * The current implementation is 1bpp RGB, with 16 pixels per SRAM word
 * Bottom 16 SRAM data bits [16; 0] are red, bit[15] leftmost
 * Next 16 SRAM data bits [16; 16] are green, bit[31] leftmost
 * Top 16 SRAM data bits [16; 132] are blue, bit[47] leftmost
 *
 */
/*a Includes */
include "apb::csr.h"
include "video::video.h"
include "apb::csr_targets.h"
include "std::srams.h"
include "video::framebuffer_modules.h"

/*a Types */
/*t t_csr_address
 *
 * CSR address decode for the framebuffer module
 */
typedef enum[4] {
    csr_address_base_address    = 0,
    csr_address_words_per_line  = 1,
} t_csr_address;

/*t t_pixel_combs 
 *
 * Combinatorial decode of the pixel_state, to determine the next
 * state
 */
typedef struct {
    bit[8] red                       "Red pixel data to be presented on the video output bus";
    bit[8] green                     "Green pixel data to be presented on the video output bus";
    bit[8] blue                      "Blue pixel data to be presented on the video output bus";
    bit[5] next_num_valid            "Number of pixels valid in the shift register after shifting or clearing at end of line";
    bit[14] sram_address_next_line   "SRAM address of the start of the next line; this is one line on from the current SRAM line start address";
    bit load_shift_register          "Asserted if the shift register is to be loaded from the data buffer";
    bit sram_request                 "Asserted if the SRAM should be read, as the data buffer is empty and data will be needed";
} t_pixel_combs;

/*t t_pixel_shift_register
 *
 * Pixel shift register contents - used for the data buffer and the shift register itself
 */
typedef struct {
    bit[16] red    "Red pixel data";
    bit[16] green  "Green pixel data";
    bit[16] blue   "Blue pixel data";
} t_pixel_shift_register;

/*t t_pixel_state
 *
 * State of the pixel logic; SRAM addresses, data buffer, shift register, and pixel data for output
 */
typedef struct {
    bit[5] num_valid                   "Number of bits valid in the shift register, from 0 to 16";
    bit[14] sram_address               "SRAM address of the next pixel data to be read";
    bit[14] sram_address_line_start    "SRAM address of the start of the current line";
    bit data_buffer_full               "Asserted if the data buffer is full";
    bit load_data_buffer               "Asserted if the SRAM read data is valid and should be loaded into the data buffer";
    t_pixel_shift_register shift       "Pixel shift register contents";
    t_pixel_shift_register data_buffer "Pixel data buffer contents";
    bit[8] red                         "Red pixel data for the @a video_bus";
    bit[8] green                       "Green pixel data for the @a video_bus";
    bit[8] blue                        "Blue pixel data for the @a video_bus";
} t_pixel_state;

/*t t_sram_state
 *
 * State in the SRAM clock domain - a buffer of the write request, to guarantee timing
*/
typedef struct {
    t_sram_access_req write_request "Write request to perform to the SRAM";
} t_sram_state;

/*t t_csrs
 *
 * Control and status register contents
 */
typedef struct {
    bit[16] sram_base_address     "Base address in SRAM of the framebuffer";
    bit[16] sram_words_per_line   "SRAM words per line used for pixel data";
    bit     down_sample_x         "Asserted if the pixel data should be down-samples by a factor of 2 (perhaps should be the 'output data mode')";
} t_csrs;

/*a Module
 */
module framebuffer( clock csr_clk "Clock for CSR reads/writes",
                    clock sram_clk  "SRAM write clock, with frame buffer data",
                    clock video_clk "Video clock, used to generate vsync, hsync, data out, etc",
                    input bit reset_n,
                    input t_sram_access_req display_sram_write,
                    output t_video_bus video_bus,
                    input t_csr_request csr_request,
                    output t_csr_response csr_response,
                    input bit[16]         csr_select
    )
"""
This is a module that takes SRAM writes into a
framebuffer, and includes a mapping to a dual-port SRAM (write on
one side, read on the other), where the video side drives out
vsync, hsync, data enable and pixel data.

The video side is asynchronous to the SRAM write side.

Video timing is handled by a @a framebuffer_timing module, which
generates the synchronization signals and display enable. This module
must be configure correctly for the display size and porches.

The video output start at a programmable base address in SRAM;
moving down a line adds a programmable amount to the address in
SRAM.

The module generates output pixel data from a shift register and a
data buffer that fill from an internal dual-port SRAM, using the video
timing.

The SRAM is filled with SRAM write requests, using a different clock
to the video generation.

The current implementation is 1bpp RGB, with 16 pixels per SRAM word
Bottom 16 SRAM data bits [16; 0] are red, bit[15] leftmost
Next 16 SRAM data bits [16; 16] are green, bit[31] leftmost
Top 16 SRAM data bits [16; 132] are blue, bit[47] leftmost

"""
{
    /*b State etc in CSR domain */
    default reset active_low reset_n;
    default clock csr_clk;
    clocked t_csrs csrs = {*=0,
                           down_sample_x=1,
                           sram_words_per_line=40 } "Control/status registers local to this module";
    net t_csr_response     csr_response_timing "Pipelined CSR response interface to control the module";
    net t_csr_response     csr_response_local  "Pipelined CSR response interface to control the module";
    net t_csr_access       csr_access          "CSR access for this module";
    comb t_csr_access_data csr_read_data       "CSR read data from this module";

    /*b State in SRAM domain */
    default reset active_low reset_n;
    default clock sram_clk;
    clocked t_sram_state    sram_state={*=0}   "State in the SRAM clock domain - the SRAM write to be performed";

    /*b State in video domain */
    default reset active_low reset_n;
    default clock video_clk;
    net t_video_timing video_timing             "Video timing syncs and controls";
    clocked t_pixel_state pixel_state={*=0}     "Pixel state, in the video clock domain, to generate the pixel data out";
    comb    t_pixel_combs pixel_combs           "Combinatorial decode of the pixel state";
    net bit[48] pixel_read_data                 "Data read from the framebuffer; currently always intepreted as bundle(16 blue, 16 green, 16 red)";

    /*b Pixel data buffer, shift register, and sram request */
    pixel_data_logic """
    The framebuffer timing is handled by a submodule; this generates
    sync and other timing signals.

    The pixel data buffer is cleared after the display portion of a
    scanline, and loaded for scanlines that are being displayed
    whenever it is empty.

    The pixel data shift register is copied from the pixel data buffer
    when it empties, and shifts down when pixels are to be displayed.

    The pixel data buffer is loaded from an SRAM, which returns data
    in the cycle after request. Hence the SRAM is read only when the
    pixel data buffer is empty _and_ the SRAM is not being read; this
    requires a minimum back porch time of about 3 clock ticks, and a
    maximum data consumption rate of one SRAM word every 3 clock
    ticks. Faster than this and the mechanism here does not keep
    up. This is not an issue currently as the maximum data consumption
    rate is with down-samping by a factor of 2 - hence 8 ticks between
    shift register emptying.
    """: {
        /*b Framebuffer timing module */
        framebuffer_timing ftiming( csr_clk <- csr_clk,
                                    video_clk <- video_clk,
                                    reset_n <= reset_n,
                                    video_timing => video_timing,
                                    csr_request <= csr_request,
                                    csr_response => csr_response_timing,
                                    csr_select <= bundle(csr_select[15;1], 1b0) );

        /*b Pixel combinatorials */
        pixel_combs.next_num_valid = pixel_state.num_valid - 1;
        if (csrs.down_sample_x) {
            pixel_combs.next_num_valid = pixel_state.num_valid - 2;
        }
        if (pixel_state.num_valid==0) {
            pixel_combs.next_num_valid = 0;
        }
        if (!video_timing.will_display_enable) {
            pixel_combs.next_num_valid = pixel_state.num_valid;
        }

        pixel_combs.sram_address_next_line  = pixel_state.sram_address_line_start + csrs.sram_words_per_line[14;0];
        pixel_combs.load_shift_register     = (pixel_state.data_buffer_full && (pixel_combs.next_num_valid==0));
        pixel_combs.sram_request            = (video_timing.v_displaying &&
                                               !(pixel_state.data_buffer_full || pixel_state.load_data_buffer) );

        pixel_combs.red   = 0;
        pixel_combs.green = 0;
        pixel_combs.blue  = 0;
        if (pixel_state.shift.red[15])   { pixel_combs.red   = -1; }
        if (pixel_state.shift.green[15]) { pixel_combs.green = -1; }
        if (pixel_state.shift.blue[15])  { pixel_combs.blue  = -1; }

        /*b Pixel state */
        pixel_state.load_data_buffer <= pixel_combs.sram_request;
        if (video_timing.will_display_enable) {
            pixel_state.shift.red[15;1]   <= pixel_state.shift.red[15;0];
            pixel_state.shift.green[15;1] <= pixel_state.shift.green[15;0];
            pixel_state.shift.blue[15;1]  <= pixel_state.shift.blue[15;0];

            if (csrs.down_sample_x) {
                pixel_state.shift.red  [14;2] <= pixel_state.shift.red  [14;0];
                pixel_state.shift.green[14;2] <= pixel_state.shift.green[14;0];
                pixel_state.shift.blue [14;2] <= pixel_state.shift.blue [14;0];
            }
            pixel_state.num_valid <= pixel_combs.next_num_valid;

            pixel_state.red   <= pixel_combs.red;
            pixel_state.green <= pixel_combs.green;
            pixel_state.blue  <= pixel_combs.blue;
        }
        if (pixel_combs.load_shift_register) {
            pixel_state.shift     <= pixel_state.data_buffer;
            pixel_state.data_buffer_full <= 0;            
            pixel_state.num_valid <= 16;
        }
        if (pixel_state.load_data_buffer) {
            pixel_state.data_buffer.red   <= pixel_read_data[16; 0];
            pixel_state.data_buffer.green <= pixel_read_data[16;16];
            pixel_state.data_buffer.blue  <= pixel_read_data[16;32];
            pixel_state.data_buffer_full <= 1;
            pixel_state.sram_address <= pixel_state.sram_address+1;
        }
        if (video_timing.will_h_sync) {
            pixel_state.data_buffer_full <= 0;            
            pixel_state.num_valid <= 0;
            if (video_timing.v_displaying) {
                pixel_state.sram_address            <= pixel_combs.sram_address_next_line;
                pixel_state.sram_address_line_start <= pixel_combs.sram_address_next_line;
            }
            if (video_timing.v_sync) {
                pixel_state.sram_address            <= csrs.sram_base_address[14;0];
                pixel_state.sram_address_line_start <= csrs.sram_base_address[14;0];
            }
        }
        /*b All done */
    }

    /*b Video bus and CSR response out */
    video_bus_out """
    The CSR responses can be combined with wire-OR; since these are
    lightweight modules there is no need to register the response for
    timing purposes.

    The video output signals come in part from the pixel state and
    from the framebuffer timing module.
    """ : {
        csr_response  = csr_response_timing;
        csr_response |= csr_response_local;

        video_bus.vsync = video_timing.v_sync;
        video_bus.hsync = video_timing.h_sync;
        video_bus.vs    = video_timing.vs;
        video_bus.hs    = video_timing.hs;
        video_bus.display_enable = video_timing.display_enable;
        video_bus.red   = pixel_state.red;
        video_bus.green = pixel_state.green;
        video_bus.blue  = pixel_state.blue;
    }
    
    /*b SRAM write and SRAM instance */
    sram_write_logic """
    Take the SRAM write bus, register it, then write in the data
    """: {
        sram_state.write_request.valid <= 0;
        if (display_sram_write.valid) {
            sram_state.write_request <= display_sram_write;
        }

        se_sram_mrw_2_16384x48 display(sram_clock_0     <- sram_clk,
                                       select_0         <= sram_state.write_request.valid,
                                       read_not_write_0 <= 0,
                                       address_0        <= sram_state.write_request.address[14;0],
                                       write_data_0     <= sram_state.write_request.write_data[48;0],
                                       // data_out_0 =>
                                       
                                       sram_clock_1     <- video_clk,
                                       select_1         <= pixel_combs.sram_request,
                                       read_not_write_1 <= 1,
                                       address_1        <= pixel_state.sram_address[14;0],
                                       write_data_1     <= 0,
                                       data_out_1       => pixel_read_data );
    }

    /*b CSR interface */
    csr_interface_logic """
    Basic read-write control status registers, using a CSR target
    interface and CSR access.
    """: {
        csr_target_csr csri( clk <- csr_clk,
                             reset_n <= reset_n,
                             csr_request  <= csr_request,
                             csr_response => csr_response_local,
                             csr_access   => csr_access,
                             csr_access_data <= csr_read_data,
                             csr_select <= bundle(csr_select[15;1], 1b1) );
        csrs <= csrs;
        csr_read_data = 0;
        part_switch (csr_access.address[4;0]) {
        case csr_address_base_address: {
            csr_read_data = bundle(16b0, csrs.sram_base_address);
            if (csr_access.valid && !csr_access.read_not_write) {
                csrs.sram_base_address   <= csr_access.data[16;0]; }
        }
        case csr_address_words_per_line: {
            csr_read_data = bundle(15b0, csrs.down_sample_x, csrs.sram_words_per_line);
            if (csr_access.valid && !csr_access.read_not_write) {
                csrs.down_sample_x         <= csr_access.data[16];
                csrs.sram_words_per_line   <= csr_access.data[16;0]; }
        }
        }

    }

    /*b All done */
}
